`ifndef DEFINE__SV
`define DEFINE__SV

//`define CALLBACK
//`define BLUEPRINT

`endif
