
`include "bp_bfm.sv"

module top;


bp_bfm bfm();





endmodule
